# ====================================================================
#
#      dharma_eth_drivers.cdl
#
#      Ethernet drivers - platform dependent support for Dharma
#                         family of development boards
#
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      toddm
# Original data:  toddm
# Contributors:
# Date:           2001-09-11
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ARM_DHARMA {
    display       "Dharma Orinoco driver"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_ARM_EDB7XXX

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH1
    include_dir   .
    include_files ; # none _exported_ whatsoever
    description   "Ethernet driver for Dharma Orinoco PC card."
#    compile       -library=libextras.a if_orinoco.c hcf.c hcfio.c
    compile       -library=libextras.a if_pc_orinoco.c hcf.c hcfio.c

    cdl_option CYGDAT_ARM_DHARMA_SET_SSID {
	display "Set the desired SSID (network name)"
	flavor  data
	default_value {"\"Todd\""}
	description "The SSID is the name of the network you with to connect to.
	NULL means to connect to any available network."
    }

    cdl_option CYGDAT_ARM_DHARMA_SET_CHANNEL {
	display "Set the channel to use"
	flavor data
	default_value {"10"}
	description "This is the channel that the driver will use to communicate."
    }

    cdl_component CYGPKG_DEVS_ETH_ARM_DHARMA_OPTIONS {
        display "Dharma Orinoco driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_ARM_DHARMA_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Dharma Orinoco driver package.
                These flags are used in addition
                to the set of global flags."
        }

	cdl_option CYGPKG_DEVS_ETH_ARM_DHARMA_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the driver. These flags are removed from
                the set of global flags if present."
        }
    }
}

