#====================================================================
#
#      flash_dharma.cdl
#
#      FLASH memory - Hardware support on IObjects dharma eval board
#
#====================================================================

cdl_package CYGPKG_DEVS_FLASH_DHARMA {
    display       "IObjects Dharma FLASH memory support"
    description   "FLASH memory device support for IObjects Dharma"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires	  CYGPKG_HAL_ARM_EDB7XXX
    implements    CYGHWR_IO_FLASH_DEVICE
    implements    CYGHWR_IO_FLASH_DEVICE_NOT_IN_RAM

    compile       dharma_flash.c dharma.c

    include_dir   cyg/io

    cdl_component CYGPKG_DEVS_FLASH_DHARMA_OPTIONS {
        display   "Flash configuration options"
        flavor    none
        no_define
        parent    CYGPKG_DEVS_FLASH_DHARMA
        
        cdl_option CYGDAT_DEVS_FLASH_DHARMA_DEVICE_SIZE {
            display     "Size of the J3 (strata) flash part being used in Mb"
            flavor      data
            default_value   128
            legal_values    128 32
            description "
              The size of the J3 part being used in Mb."
        }
        cdl_option CYGNUM_DEVS_FLASH_DHARMA_NUM_DEVICES {
            display     "Number of J3 devices"
            flavor      data
            default_value   2
            legal_values    1 2
            description "
                The number of J3 devices being used. 1 for 16-bit configurations, 2 for 32-bit."
        }
    }

    make -priority 1 {
        flash_erase_block.o: $(REPOSITORY)/$(PACKAGE)/src/flash_erase_block.c \
                             $(REPOSITORY)/$(PACKAGE)/src/dharma.h
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_erase_block.c
        echo " .globl flash_erase_block_end" >>flash_erase_block.s
        echo "flash_erase_block_end:" >>flash_erase_block.s
        $(CC) -c -o flash_erase_block.o flash_erase_block.s
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_erase_block.o
    }
    make -priority 1 {
        flash_program_buf.o: $(REPOSITORY)/$(PACKAGE)/src/flash_program_buf.c \
                             $(REPOSITORY)/$(PACKAGE)/src/dharma.h
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_program_buf.c
        echo " .globl flash_program_buf_end" >>flash_program_buf.s
        echo "flash_program_buf_end:" >>flash_program_buf.s
        $(CC) -c -o flash_program_buf.o flash_program_buf.s
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_program_buf.o
    }
    make -priority 1 {
        flash_query.o: $(REPOSITORY)/$(PACKAGE)/src/flash_query.c \
                             $(REPOSITORY)/$(PACKAGE)/src/dharma.h
        $(CC) -S $(INCLUDE_PATH) $(CFLAGS) -g0 -fno-function-sections $(REPOSITORY)/$(PACKAGE)/src/flash_query.c
        echo " .globl flash_query_end" >>flash_query.s
        echo "flash_query_end:" >>flash_query.s
        $(CC) -c -o flash_query.o flash_query.s
        $(AR) rcs $(PREFIX)/lib/libtarget.a flash_query.o
    }

}
