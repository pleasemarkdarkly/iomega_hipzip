# ====================================================================
#
#      edb7xxx_eth_drivers.cdl
#
#      Ethernet drivers - platform dependent support for Cirrus Logic
#                         EDB7xxx family of development boards
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, jskov
# Date:           2000-01-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ARM_EDB7XXX {
    display       "Cirrus Logic ethernet driver for EP7xxx boards"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_ARM_EDB7XXX

    include_dir   cyg/io

    description   "Ethernet driver for Cirrus Logic EP7xxx based
                  development boards."

    # FIXME: This really belongs in the CL CS8900A package
    cdl_interface CYGINT_DEVS_ETH_CL_CS8900A_REQUIRED {
        display   "Cirrus Logic CS8900A ethernet driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_CL_CS8900A_INL <cyg/io/devs_eth_arm_edb7xxx.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_CL_CS8900A_CFG <pkgconf/devs_eth_arm_edb7xxx.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }

    cdl_component CYGPKG_DEVS_ETH_ARM_EDB7XXX_ETH0 {
        display       "EDB7XXX ethernet port driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the ethernet device driver for the
            EDB7XXX port."

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH0
        implements CYGINT_DEVS_ETH_CL_CS8900A_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_ARM_EDB7XXX_ETH0_NAME {
            display       "Device name for the ETH0 ethernet driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device."
        }

        cdl_option CYGDAT_DEVS_ETH_ARM_EDB7XXX_ETH0_BASE_ADDRESS {
            display       "Set the controller base address"
            flavor        data
            default_value { CYGHWR_HAL_ARM_EDB7XXX_BOARD_VARIANT == "DHARMA_V2" ? 0xf0000000 :
                            0x20000000 }
            description   "This option sets the base address for the
            ethernet controller. This is useful for hardware spins that
            put the same device on a different chip select."
        }
        cdl_component CYGSEM_DEVS_ETH_ARM_EDB7XXX_ETH0_SET_ESA {
            display       "Set the ethernet station address"
            flavor        bool
            calculated    0
            description   "Enabling this option will allow the ethernet
            station address to be forced to the value set by the
            configuration.  This may be required if the hardware does
            not include a serial EEPROM for the ESA."
            
            cdl_option CYGDAT_DEVS_ETH_ARM_EDB7XXX_ETH0_ESA {
                display       "The ethernet station address"
                flavor        data
                default_value {"{0x08, 0x88, 0x12, 0x34, 0x56, 0x78}"}
                description   "The ethernet station address"
            }
        }
    }

}

